/*
 *  
 *  Copyright(C) 2018 Gerald Coe, Devantech Ltd <gerry@devantech.co.uk>
 * 
 *  Permission to use, copy, modify, and/or distribute this software for any purpose with or
 *  without fee is hereby granted, provided that the above copyright notice and 
 *  this permission notice appear in all copies.
 * 
 *  THE SOFTWARE IS PROVIDED "AS IS" AND THE AUTHOR DISCLAIMS ALL WARRANTIES WITH REGARD TO
 *  THIS SOFTWARE INCLUDING ALL IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS. 
 *  IN NO EVENT SHALL THE AUTHOR BE LIABLE FOR ANY SPECIAL, DIRECT, INDIRECT, OR CONSEQUENTIAL 
 *  DAMAGES OR ANY DAMAGES WHATSOEVER RESULTING FROM LOSS OF USE, DATA OR PROFITS, WHETHER IN
 *  AN ACTION OF CONTRACT, NEGLIGENCE OR OTHER TORTIOUS ACTION, ARISING OUT OF OR IN 
 *  CONNECTION WITH THE USE OR PERFORMANCE OF THIS SOFTWARE.
 * 
 */
 


module LedStrip (
	input clk12MHz,
	input [7:0] RedPWM,
	input [7:0] GreenPWM,
	input [7:0] BluePWM,
	output reg Red,
	output reg Green,
	output reg Blue 
	);

	reg [7:0] timer;
	
	always @ (posedge clk12MHz) begin
		timer <= timer+1;
		if(RedPWM==timer) Red <= 1'b0;
		else if(timer==8'b0) Red <= 1'b1;
		else Red <= Red;

		if(GreenPWM==timer) Green <= 1'b0;
		else if(timer==8'b0) Green <= 1'b1;
		else Green <= Green;

		if(BluePWM==timer) Blue <= 1'b0;
		else if(timer==8'b0) Blue <= 1'b1;
		else Blue <= Blue;
	end

endmodule



